----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:04:10 05/27/2021 
-- Design Name: 
-- Module Name:    vga1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------

LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
USE ieee.std_logic_signed.all ;
USE ieee.std_logic_arith.all ;
USE ieee.std_logic_unsigned.all;
entity ee240_vgadriver is
		port (
			nreset: in std_logic;
			board_clk: in std_logic;
			vsync: out std_logic;
			hsync: out std_logic;
			red: out std_logic_vector(2 downto 0);
			green: out std_logic_vector(2 downto 0);
			blue: out std_logic_vector(1 downto 0)
		);
end;

architecture arch_vga_driver of ee240_vgadriver is

component freq_divider 
	port(
	board_clock : in std_logic;
	reset: in std_logic;
	divided_clock: out std_logic
	);
end component;

component horizontal_sync_generator 
	port(
		clock: in std_logic;
		reset: in std_logic;
		hsync: out std_logic;
		communicate_vsync: out std_logic;
		display_enable_H: out std_logic
	);
end component;

component vertical_sync_generator
	port(
		clock: in std_logic;
		reset: in std_logic;
		vsync: out std_logic;
		communicate_color_gen: out std_logic;
		display_enable_V: out std_logic
	);
end component;

component color_generator 
	port(
	clock: in std_logic;
	reset: in std_logic;
	colors: out std_logic_vector (7 downto 0)
	);
end component;

signal clock25MHz : std_logic; --this signal stores the processed clock cycle which is 25 MHz from 100 MHz clock
signal horizontal_sync: std_logic; --this signal stores the horizontal signal described in lab guide
signal vertical_sync: std_logic; --this signal stores the vertical signal described in lab guide
signal horizontal_gen_period_complete: std_logic; --this signal an impulse which becomes 1 when the period of the horizontal signal is completed and then becomes immediately 0
--one of the overall horizontal signal corresponds to one clock cycle for  the vertical generator, that's why horizontal period complete signal is used for the clock for the vertical sync. gen
signal vertical_gen_period_complete: std_logic; --this signal an impulse which becomes 1 when the period of the vertical signal is completed and then becomes immediately 0
--one of the overall vertical signal corresponds to the one frame on a screen, so after completing this period frame normally changes, I connected this impulse signal to the reset of the color in order to reset it before another frame comes in
signal horizontal_sync_color_enable: std_logic;
--it is 1 when T_disp is 1 for the horizontal sync signal (which allows screen to display correct color in right place)
signal vertical_sync_color_enable: std_logic;
--it is 1 when T_disp is 1 for the horizontal sync signal (which allows screen to display correct color in right place)
signal vertical_and_horizontal_sync_to_color_gen: std_logic;
--this signal represents the reset signal of the color gen : which consists of the not (T_disp of the hsync and vsync) with the period done signal of  vsync
signal resulting_colors: std_logic_vector(7 downto 0);
--stores the color bits generated by the color generator will be intermediate signal between the output and the generator (just created to make more obvious of main module)
begin

 f1: freq_divider port map(board_clk,nreset,clock25MHz);
--freq divider takes the  board clock (100MHz => )and reset signal and generates 25MHz clock 
 f2: horizontal_sync_generator port map (clock25MHz,nreset,horizontal_sync,horizontal_gen_period_complete,horizontal_sync_color_enable);
 --takes the 25MHz clock and generates corresponding signals indicated at the above
 f3: vertical_sync_generator port map (horizontal_gen_period_complete,nreset,vertical_sync, vertical_gen_period_complete,vertical_sync_color_enable);
 --takes the horizontal period done signal as clock and generates corresponding singals indicated at the above
 vertical_and_horizontal_sync_to_color_gen <= not (horizontal_sync_color_enable and vertical_sync_color_enable) or vertical_gen_period_complete;
 -- color signal should be set whenever one of the T_disps of the sync generators is 0 or period is done by vsync (period os vysync is not necessary if frame doesn't changes)
 f4: color_generator port map(clock25MHz, vertical_and_horizontal_sync_to_color_gen,resulting_colors);
 --generates color signal with 25MHz bit clock and according to the respective reset signal 
 
 --assigning generated signals to th outputs starts here:
 HSYNC <= horizontal_sync;
 VSYNC <= vertical_sync;
 red <= resulting_colors (7 downto 5);
 green <= resulting_colors (4 downto 2);
 blue <= resulting_colors (1 downto 0);
 --ends here:
 
-- nreset comes from BTNS (Push-Button Switch) 
-- board_clk comes from the 100 MHz board clock
--vsync is connected to VGA-VSYNC#
--hsync is connected to VGA-HSYNC#
--red(0) is connected to VGA-RED0
--red(1) is connected to VGA-RED1
--red(2) is connected to VGA-RED2
--green(0) is connected to VGA-GRN0
--green(1) is connected to VGA-GRN1
--green(2) is connected to VGA-GRN2
--blue(0) is connected to VGA-BLU1
--blue(1) is connected to VGA-BLU2
end arch_vga_driver;
